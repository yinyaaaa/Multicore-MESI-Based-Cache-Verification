`define INST_TOP_CORE inst_cache_lv1_multicore
`define NUM_CORE 4
`define DATA_ADDR_START 32'h4000_0000