//=====================================================================
// Project: 4 core MESI cache design
// File Name: read_miss_icache.sv
// Description: Test for read-miss to I-cache
// Designers: Venky & Suru
//=====================================================================

class lru extends base_test;

    //component macro
    `uvm_component_utils(lru)

    //Constructor
    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction : new

    //UVM build phase
    function void build_phase(uvm_phase phase);
        uvm_config_wrapper::set(this, "tb.vsequencer.run_phase", "default_sequence", lru_seq::type_id::get());
        super.build_phase(phase);
    endfunction : build_phase

    //UVM run phase()
    task run_phase(uvm_phase phase);
        `uvm_info(get_type_name(), "Executing lru test" , UVM_LOW)
    endtask: run_phase

endclass : lru


// Sequence for a read-miss on I-cache
class lru_seq extends base_vseq;
    //object macro
    `uvm_object_utils(lru_seq)

    cpu_transaction_c trans;

    //constructor
    function new (string name="lru_seq");
        super.new(name);
    endfunction : new

    virtual task body();
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == WRITE_REQ; address == 32'h5000_AAAA; data == 32'h0000_0001;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == WRITE_REQ; address == 32'h6000_AAAA; data == 32'h0000_0002;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == WRITE_REQ; address == 32'h7000_AAAA; data == 32'h0000_0003;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == WRITE_REQ; address == 32'h8000_AAAA; data == 32'h0000_0004;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == WRITE_REQ; address == 32'h9000_AAAA; data == 32'h0000_0005;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == WRITE_REQ; address == 32'ha000_AAAA; data == 32'h0000_0006;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == WRITE_REQ; address == 32'hb000_AAAA; data == 32'h0000_0007;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == WRITE_REQ; address == 32'hc000_AAAA; data == 32'h0000_0008;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == READ_REQ; address == 32'h5000_AAAA;}) 
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == READ_REQ; address == 32'h6000_AAAA;}) 
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == READ_REQ; address == 32'h7000_AAAA;}) 
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0],{request_type == READ_REQ; address == 32'h8000_AAAA;}) 

    endtask

endclass : lru_seq
